//MIT License
//
//Copyright (c) 2024 Yuri Korotaev
//
//Permission is hereby granted, free of charge, to any person obtaining a copy
//of this software and associated documentation files (the "Software"), to deal
//in the Software without restriction, including without limitation the rights
//to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
//copies of the Software, and to permit persons to whom the Software is
//furnished to do so, subject to the following conditions:
//
//The above copyright notice and this permission notice shall be included in all
//copies or substantial portions of the Software.
//
//THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
//IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
//FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
//AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
//LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
//OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
//SOFTWARE.

module APUF_Cyclone4

# (parameter line_length = 3)

(
    input clk,
    input [line_length - 1 :0] challenge,

    output response

);

wire delay_line_out_1;
wire delay_line_out_2;


delay_line delay_line(
    .clk(clk),
    .challenge(challenge),
    .line_out_1(delay_line_out_1),
    .line_out_2(delay_line_out_2)
);

dff dff(
    .clk(delay_line_out_2),
    .d(delay_line_out_1),
    .q(response)
);

endmodule